`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/05/12 15:30:21
// Design Name: 
// Module Name: Sbox
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sbox(in,id,out);
    input [5:0]in;
    input [3:0]id;
    output [3:0]out;
    assign out=SBOX(in,id);
    function [4:1] SBOX(input [6:1] B, input reg [4:0] s_table_id);

    reg [2:1] i;

    reg [4:1] j;

    reg [3:0] S1[3:0][15:0];

    reg [3:0] S2[3:0][15:0];

    reg [3:0] S3[3:0][15:0];

    reg [3:0] S4[3:0][15:0];

    reg [3:0] S5[3:0][15:0];

    reg [3:0] S6[3:0][15:0];

    reg [3:0] S7[3:0][15:0];

    reg [3:0] S8[3:0][15:0];

    begin

			S1[0][0] = 14;

			S1[0][1] = 4;

			S1[0][2] = 13;

			S1[0][3] = 1;

			S1[0][4] = 2;

			S1[0][5] = 15;

			S1[0][6] = 11;

			S1[0][7] = 8;

			S1[0][8] = 3;

			S1[0][9] = 10;

			S1[0][10] = 6;

			S1[0][11] = 12;

			S1[0][12] = 5;

			S1[0][13] = 9;

			S1[0][14] = 0;

			S1[0][15] = 7;

			S1[1][0] = 0;

			S1[1][1] = 15;

			S1[1][2] = 7;

			S1[1][3] = 4;

			S1[1][4] = 14;

			S1[1][5] = 2;

			S1[1][6] = 13;

			S1[1][7] = 1;

			S1[1][8] = 10;

			S1[1][9] = 6;

			S1[1][10] = 12;

			S1[1][11] = 11;

			S1[1][12] = 9;

			S1[1][13] = 5;

			S1[1][14] = 3;

			S1[1][15] = 8;

			S1[2][0] = 4;

			S1[2][1] = 1;

			S1[2][2] = 14;

			S1[2][3] = 8;

			S1[2][4] = 13;

			S1[2][5] = 6;

			S1[2][6] = 2;

			S1[2][7] = 11;

			S1[2][8] = 15;

			S1[2][9] = 12;

			S1[2][10] = 9;

			S1[2][11] = 7;

			S1[2][12] = 3;

			S1[2][13] = 10;

			S1[2][14] = 5;

			S1[2][15] = 0;

			S1[3][0] = 15;

			S1[3][1] = 12;

			S1[3][2] = 8;

			S1[3][3] = 2;

			S1[3][4] = 4;

			S1[3][5] = 9;

			S1[3][6] = 1;

			S1[3][7] = 7;

			S1[3][8] = 5;

			S1[3][9] = 11;

			S1[3][10] = 3;

			S1[3][11] = 14;

			S1[3][12] = 10;

			S1[3][13] = 0;

			S1[3][14] = 6;

			S1[3][15] = 13;

			S2[0][0] = 15;

			S2[0][1] = 1;

			S2[0][2] = 8;

			S2[0][3] = 14;

			S2[0][4] = 6;

			S2[0][5] = 11;

			S2[0][6] = 3;

			S2[0][7] = 4;

			S2[0][8] = 9;

			S2[0][9] = 7;

			S2[0][10] = 2;

			S2[0][11] = 13;

			S2[0][12] = 12;

			S2[0][13] = 0;

			S2[0][14] = 5;

			S2[0][15] = 10;

			S2[1][0] = 3;

			S2[1][1] = 13;

			S2[1][2] = 4;

			S2[1][3] = 7;

			S2[1][4] = 15;

			S2[1][5] = 2;

			S2[1][6] = 8;

			S2[1][7] = 14;

			S2[1][8] = 12;

			S2[1][9] = 0;

			S2[1][10] = 1;

			S2[1][11] = 10;

			S2[1][12] = 6;

			S2[1][13] = 9;

			S2[1][14] = 11;

			S2[1][15] = 5;

			S2[2][0] = 0;

			S2[2][1] = 14;

			S2[2][2] = 7;

			S2[2][3] = 11;

			S2[2][4] = 10;

			S2[2][5] = 4;

			S2[2][6] = 13;

			S2[2][7] = 1;

			S2[2][8] = 5;

			S2[2][9] = 8;

			S2[2][10] = 12;

			S2[2][11] = 6;

			S2[2][12] = 9;

			S2[2][13] = 3;

			S2[2][14] = 2;

			S2[2][15] = 15;

			S2[3][0] = 13;

			S2[3][1] = 8;

			S2[3][2] = 10;

			S2[3][3] = 1;

			S2[3][4] = 3;

			S2[3][5] = 15;

			S2[3][6] = 4;

			S2[3][7] = 2;

			S2[3][8] = 11;

			S2[3][9] = 6;

			S2[3][10] = 7;

			S2[3][11] = 12;

			S2[3][12] = 0;

			S2[3][13] = 5;

			S2[3][14] = 14;

			S2[3][15] = 9;

			S3[0][0] = 10;

			S3[0][1] = 0;

			S3[0][2] = 9;

			S3[0][3] = 14;

			S3[0][4] = 6;

			S3[0][5] = 3;

			S3[0][6] = 15;

			S3[0][7] = 5;

			S3[0][8] = 1;

			S3[0][9] = 13;

			S3[0][10] = 12;

			S3[0][11] = 7;

			S3[0][12] = 11;

			S3[0][13] = 4;

			S3[0][14] = 2;

			S3[0][15] = 8;

			S3[1][0] = 13;

			S3[1][1] = 7;

			S3[1][2] = 0;

			S3[1][3] = 9;

			S3[1][4] = 3;

			S3[1][5] = 4;

			S3[1][6] = 6;

			S3[1][7] = 10;

			S3[1][8] = 2;

			S3[1][9] = 8;

			S3[1][10] = 5;

			S3[1][11] = 14;

			S3[1][12] = 12;

			S3[1][13] = 11;

			S3[1][14] = 15;

			S3[1][15] = 1;

			S3[2][0] = 13;

			S3[2][1] = 6;

			S3[2][2] = 4;

			S3[2][3] = 9;

			S3[2][4] = 8;

			S3[2][5] = 15;

			S3[2][6] = 3;

			S3[2][7] = 0;

			S3[2][8] = 11;

			S3[2][9] = 1;

			S3[2][10] = 2;

			S3[2][11] = 12;

			S3[2][12] = 5;

			S3[2][13] = 10;

			S3[2][14] = 14;

			S3[2][15] = 7;

			S3[3][0] = 1;

			S3[3][1] = 10;

			S3[3][2] = 13;

			S3[3][3] = 0;

			S3[3][4] = 6;

			S3[3][5] = 9;

			S3[3][6] = 8;

			S3[3][7] = 7;

			S3[3][8] = 4;

			S3[3][9] = 15;

			S3[3][10] = 14;

			S3[3][11] = 3;

			S3[3][12] = 11;

			S3[3][13] = 5;

			S3[3][14] = 2;

			S3[3][15] = 12;

			S4[0][0] = 7;

			S4[0][1] = 13;

			S4[0][2] = 14;

			S4[0][3] = 3;

			S4[0][4] = 0;

			S4[0][5] = 6;

			S4[0][6] = 9;

			S4[0][7] = 10;

			S4[0][8] = 1;

			S4[0][9] = 2;

			S4[0][10] = 8;

			S4[0][11] = 5;

			S4[0][12] = 11;

			S4[0][13] = 12;

			S4[0][14] = 4;

			S4[0][15] = 15;

			S4[1][0] = 13;

			S4[1][1] = 8;

			S4[1][2] = 11;

			S4[1][3] = 5;

			S4[1][4] = 6;

			S4[1][5] = 15;

			S4[1][6] = 0;

			S4[1][7] = 3;

			S4[1][8] = 4;

			S4[1][9] = 7;

			S4[1][10] = 2;

			S4[1][11] = 12;

			S4[1][12] = 1;

			S4[1][13] = 10;

			S4[1][14] = 14;

			S4[1][15] = 9;

			S4[2][0] = 10;

			S4[2][1] = 6;

			S4[2][2] = 9;

			S4[2][3] = 0;

			S4[2][4] = 12;

			S4[2][5] = 11;

			S4[2][6] = 7;

			S4[2][7] = 13;

			S4[2][8] = 15;

			S4[2][9] = 1;

			S4[2][10] = 3;

			S4[2][11] = 14;

			S4[2][12] = 5;

			S4[2][13] = 2;

			S4[2][14] = 8;

			S4[2][15] = 4;

			S4[3][0] = 3;

			S4[3][1] = 15;

			S4[3][2] = 0;

			S4[3][3] = 6;

			S4[3][4] = 10;

			S4[3][5] = 1;

			S4[3][6] = 13;

			S4[3][7] = 8;

			S4[3][8] = 9;

			S4[3][9] = 4;

			S4[3][10] = 5;

			S4[3][11] = 11;

			S4[3][12] = 12;

			S4[3][13] = 7;

			S4[3][14] = 2;

			S4[3][15] = 14;

			S5[0][0] = 2;

			S5[0][1] = 12;

			S5[0][2] = 4;

			S5[0][3] = 1;

			S5[0][4] = 7;

			S5[0][5] = 10;

			S5[0][6] = 11;

			S5[0][7] = 6;

			S5[0][8] = 8;

			S5[0][9] = 5;

			S5[0][10] = 3;

			S5[0][11] = 15;

			S5[0][12] = 13;

			S5[0][13] = 0;

			S5[0][14] = 14;

			S5[0][15] = 9;

			S5[1][0] = 14;

			S5[1][1] = 11;

			S5[1][2] = 2;

			S5[1][3] = 12;

			S5[1][4] = 4;

			S5[1][5] = 7;

			S5[1][6] = 13;

			S5[1][7] = 1;

			S5[1][8] = 5;

			S5[1][9] = 0;

			S5[1][10] = 15;

			S5[1][11] = 10;

			S5[1][12] = 3;

			S5[1][13] = 9;

			S5[1][14] = 8;

			S5[1][15] = 6;

			S5[2][0] = 4;

			S5[2][1] = 2;

			S5[2][2] = 1;

			S5[2][3] = 11;

			S5[2][4] = 10;

			S5[2][5] = 13;

			S5[2][6] = 7;

			S5[2][7] = 8;

			S5[2][8] = 15;

			S5[2][9] = 9;

			S5[2][10] = 12;

			S5[2][11] = 5;

			S5[2][12] = 6;

			S5[2][13] = 3;

			S5[2][14] = 0;

			S5[2][15] = 14;

			S5[3][0] = 11;

			S5[3][1] = 8;

			S5[3][2] = 12;

			S5[3][3] = 7;

			S5[3][4] = 1;

			S5[3][5] = 14;

			S5[3][6] = 2;

			S5[3][7] = 13;

			S5[3][8] = 6;

			S5[3][9] = 15;

			S5[3][10] = 0;

			S5[3][11] = 9;

			S5[3][12] = 10;

			S5[3][13] = 4;

			S5[3][14] = 5;

			S5[3][15] = 3;

			S6[0][0] = 12;

			S6[0][1] = 1;

			S6[0][2] = 10;

			S6[0][3] = 15;

			S6[0][4] = 9;

			S6[0][5] = 2;

			S6[0][6] = 6;

			S6[0][7] = 8;

			S6[0][8] = 0;

			S6[0][9] = 13;

			S6[0][10] = 3;

			S6[0][11] = 4;

			S6[0][12] = 14;

			S6[0][13] = 7;

			S6[0][14] = 5;

			S6[0][15] = 11;

			S6[1][0] = 10;

			S6[1][1] = 15;

			S6[1][2] = 4;

			S6[1][3] = 2;

			S6[1][4] = 7;

			S6[1][5] = 12;

			S6[1][6] = 9;

			S6[1][7] = 5;

			S6[1][8] = 6;

			S6[1][9] = 1;

			S6[1][10] = 13;

			S6[1][11] = 14;

			S6[1][12] = 0;

			S6[1][13] = 11;

			S6[1][14] = 3;

			S6[1][15] = 8;

			S6[2][0] = 9;

			S6[2][1] = 14;

			S6[2][2] = 15;

			S6[2][3] = 5;

			S6[2][4] = 2;

			S6[2][5] = 8;

			S6[2][6] = 12;

			S6[2][7] = 3;

			S6[2][8] = 7;

			S6[2][9] = 0;

			S6[2][10] = 4;

			S6[2][11] = 10;

			S6[2][12] = 1;

			S6[2][13] = 13;

			S6[2][14] = 11;

			S6[2][15] = 6;

			S6[3][0] = 4;

			S6[3][1] = 3;

			S6[3][2] = 2;

			S6[3][3] = 12;

			S6[3][4] = 9;

			S6[3][5] = 5;

			S6[3][6] = 15;

			S6[3][7] = 10;

			S6[3][8] = 11;

			S6[3][9] = 14;

			S6[3][10] = 1;

			S6[3][11] = 7;

			S6[3][12] = 6;

			S6[3][13] = 0;

			S6[3][14] = 8;

			S6[3][15] = 13;

			S7[0][0] = 4;

			S7[0][1] = 11;

			S7[0][2] = 2;

			S7[0][3] = 14;

			S7[0][4] = 15;

			S7[0][5] = 0;

			S7[0][6] = 8;

			S7[0][7] = 13;

			S7[0][8] = 3;

			S7[0][9] = 12;

			S7[0][10] = 9;

			S7[0][11] = 7;

			S7[0][12] = 5;

			S7[0][13] = 10;

			S7[0][14] = 6;

			S7[0][15] = 1;

			S7[1][0] = 13;

			S7[1][1] = 0;

			S7[1][2] = 11;

			S7[1][3] = 7;

			S7[1][4] = 4;

			S7[1][5] = 9;

			S7[1][6] = 1;

			S7[1][7] = 10;

			S7[1][8] = 14;

			S7[1][9] = 3;

			S7[1][10] = 5;

			S7[1][11] = 12;

			S7[1][12] = 2;

			S7[1][13] = 15;

			S7[1][14] = 8;

			S7[1][15] = 6;

			S7[2][0] = 1;

			S7[2][1] = 4;

			S7[2][2] = 11;

			S7[2][3] = 13;

			S7[2][4] = 12;

			S7[2][5] = 3;

			S7[2][6] = 7;

			S7[2][7] = 14;

			S7[2][8] = 10;

			S7[2][9] = 15;

			S7[2][10] = 6;

			S7[2][11] = 8;

			S7[2][12] = 0;

			S7[2][13] = 5;

			S7[2][14] = 9;

			S7[2][15] = 2;

			S7[3][0] = 6;

			S7[3][1] = 11;

			S7[3][2] = 13;

			S7[3][3] = 8;

			S7[3][4] = 1;

			S7[3][5] = 4;

			S7[3][6] = 10;

			S7[3][7] = 7;

			S7[3][8] = 9;

			S7[3][9] = 5;

			S7[3][10] = 0;

			S7[3][11] = 15;

			S7[3][12] = 14;

			S7[3][13] = 2;

			S7[3][14] = 3;

			S7[3][15] = 12;

			S8[0][0] = 13;

			S8[0][1] = 2;

			S8[0][2] = 8;

			S8[0][3] = 4;

			S8[0][4] = 6;

			S8[0][5] = 15;

			S8[0][6] = 11;

			S8[0][7] = 1;

			S8[0][8] = 10;

			S8[0][9] = 9;

			S8[0][10] = 3;

			S8[0][11] = 14;

			S8[0][12] = 5;

			S8[0][13] = 0;

			S8[0][14] = 12;

			S8[0][15] = 7;

			S8[1][0] = 1;

			S8[1][1] = 15;

			S8[1][2] = 13;

			S8[1][3] = 8;

			S8[1][4] = 10;

			S8[1][5] = 3;

			S8[1][6] = 7;

			S8[1][7] = 4;

			S8[1][8] = 12;

			S8[1][9] = 5;

			S8[1][10] = 6;

			S8[1][11] = 11;

			S8[1][12] = 0;

			S8[1][13] = 14;

			S8[1][14] = 9;

			S8[1][15] = 2;

			S8[2][0] = 7;

			S8[2][1] = 11;

			S8[2][2] = 4;

			S8[2][3] = 1;

			S8[2][4] = 9;

			S8[2][5] = 12;

			S8[2][6] = 14;

			S8[2][7] = 2;

			S8[2][8] = 0;

			S8[2][9] = 6;

			S8[2][10] = 10;

			S8[2][11] = 13;

			S8[2][12] = 15;

			S8[2][13] = 3;

			S8[2][14] = 5;

			S8[2][15] = 8;

			S8[3][0] = 2;

			S8[3][1] = 1;

			S8[3][2] = 14;

			S8[3][3] = 7;

			S8[3][4] = 4;

			S8[3][5] = 10;

			S8[3][6] = 8;

			S8[3][7] = 13;

			S8[3][8] = 15;

			S8[3][9] = 12;

			S8[3][10] = 9;

			S8[3][11] = 0;

			S8[3][12] = 3;

			S8[3][13] = 5;

			S8[3][14] = 6;

			S8[3][15] = 11;

      

      i[2:1] = {B[6], B[1]};

      j[4:1] = B[5:2];

      

      case(s_table_id)

        5'b01: SBOX = S1[i][j];

        5'b10: SBOX = S2[i][j];

        5'b11: SBOX = S3[i][j];

        5'b100: SBOX = S4[i][j];

        5'b101: SBOX = S5[i][j];

        5'b110: SBOX = S6[i][j];

        5'b111: SBOX = S7[i][j];

        5'b1000: SBOX = S8[i][j];

      endcase

      

    end

  endfunction


endmodule
